import_C("json_struct.h");

signature sJSMN{
  void json_open( void );
  void json_parse(
    [out,size_is(btr)] char_t *c_path,
    [out,size_is(btr)] char_t *e_path,
    [out,size_is(btr)] char_t *f_path,
    [in] int btr );
  void json_arg( [out,size_is(btr)] struct arg *obj, [in] int btr );
};

celltype tJSMN {
  entry sJSMN eJSMN;
  attr{
    int16_t LEN = 256;
  };
  var {
    [size_is(LEN)]
      char_t  *json_str;
  };
};
