/* POSIX 用の簡単なテスト環境のコンポーネント記述を取り込む */
import( <cygwin_kernel.cdl> );

/* tTECSUnit セルタイプ (コンポーネントの型) */
celltype tTECSUnit {
	entry sTaskBody eMain;
};

/* TECSUnit セル (コンポーネント) */
cell tTECSUnit TECSUnit {
  /*----- TECSUnit test -----*/
};

/* Task セル (コンポーネント) */
cell tTask Task {
	cBody = TECSUnit.eMain;
	priority = 11;		/* この値は使われていない */
	stackSize = 4096;	/* この値は使われていない */
	taskAttribute = C_EXP( "TA_ACT");
};
