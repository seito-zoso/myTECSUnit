signature sTarget1 {
  int double([in] int arg);
};

signature sTarget2 {
  int add([in] int arg1, [in] int arg2);
};

celltype tTarget1 {
  entry sTarget1 eTarget1;
};

celltype tTarget2 {
  entry sTarget2 eTarget2;
};


cell tTarget1 Target1 {

};
cell tTarget2 Target2 {

};
