import_C("json_struct.h");

signature sJSMN{
  ER json_open( void );
  ER json_parse(
    [out,size_is(btr)] char_t *c_path,
    [out,size_is(btr)] char_t *e_path,
    [out,size_is(btr)] char_t *f_path,
    [in] int target_num,
    [in] int btr );
  ER json_arg(
    [out,size_is(btr)] struct tecsunit_obj *arguments,
    [out,size_is(btr)] struct tecsunit_obj *exp_val,
    [in] int target_num,
    [in] int btr );
};

celltype tJSMN {
  entry sJSMN eJSMN;
  attr{
    int16_t LEN = 256;
    char_t *key_cell = "cell";
    char_t *key_entry = "entry";
    char_t *key_function = "function";
    char_t *key_arg = "argument";
    char_t *key_exp = "exp_val";
  };
  var {
    [size_is(LEN)]
      char_t  *json_str;
    int pointer;
  };
};
