celltype tTECSUnit {
  [dynamic, optional]
    call sTest cUnitTest1;
  [dynamic, optional]
    call sTest cUnitTest2;
};
